package top_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import i2c_vip_pkg::*;

    `include "my_env.sv"
    `include "my_sequence.sv"
    `include "my_test.sv"

endpackage
