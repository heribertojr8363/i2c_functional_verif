package top_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import i2c_pkg::*;

    `include "../tb/my_env.sv"
    `include "../tb/my_test.sv"

endpackage
